`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:00:35 12/31/2020 
// Design Name: 
// Module Name:    vgaDisplayModule 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: call ip cores and vga to display objects
//
//////////////////////////////////////////////////////////////////////////////////
module vgaTop();


endmodule
