`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:01:48 12/31/2020 
// Design Name: 
// Module Name:    imgDisplayModule 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: call vgaTop
//
//////////////////////////////////////////////////////////////////////////////////
module imgDisplayModule();

	vgaTop vga();

endmodule
